library IEEE;
use  IEEE.STD_LOGIC_1164.all;

ENTITY CHECKER IS
PORT( PIPE1,PIPE2,PIPE3 : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
	PIPE1X, PIPE1G, PIPE2X, PIPE2G, PIPE3X, PIPE3G : OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END ENTITY CHECKER;

ARCHITECTURE BEHAV OF CHECKER IS
	SIGNAL IS_SAME : STD_LOGIC;
BEGIN
	IS_SAME <= '1' WHEN ( (PIPE1(8 DOWNTO 6) = PIPE2(2 DOWNTO 0)) OR (PIPE1(8 DOWNTO 6) = PIPE3(5 DOWNTO 3)) 
	OR (PIPE2(2 DOWNTO 0) = PIPE3(5 DOWNTO 3)) ) ELSE '0';

PIPE1X <= PIPE1(8 DOWNTO 6) WHEN IS_SAME='0' ELSE "000";
PIPE2X <= PIPE2(2 DOWNTO 0) WHEN IS_SAME='0' ELSE "010";
PIPE3X <= PIPE3(5 DOWNTO 3) WHEN IS_SAME='0' ELSE "100";

PIPE1G <= PIPE1(5 DOWNTO 3);
PIPE2G <= PIPE2(8 DOWNTO 6);
PIPE3G <= PIPE3(2 DOWNTO 0);

END ARCHITECTURE BEHAV;