library IEEE;
use  IEEE.STD_LOGIC_1164.all;

ENTITY LFSR_PLACEHOLDER IS
	PORT(	PIPE1_GAP, PIPE2_GAP, PIPE3_GAP, PIPE1_ENDX, 
		PIPE2_ENDX, PIPE3_ENDX : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)	
		
		);


END ENTITY LFSR_PLACEHOLDER;

ARCHITECTURE BEHAV OF LFSR_PLACEHOLDER IS

BEGIN
	PIPE1_GAP <= "000";
	PIPE2_GAP <= "001";
	PIPE3_GAP <= "010";

	PIPE1_ENDX <= "000";
	PIPE2_ENDX <= "001";
	PIPE3_ENDX <= "010";

END ARCHITECTURE BEHAV;