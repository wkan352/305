LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE IEEE.STD_LOGIC_UNSIGNED.all;
USE IEEE.NUMERIC_STD.ALL;

ENTITY D2_4bit IS
    PORT (
        VERT_SYNC : IN STD_LOGIC;
        SCORE_IN : IN INTEGER RANGE 0 TO 9;
        SCORE_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
        --Enable_OUT: OUT STD_LOGIC);
END ENTITY D2_4bit;

ARCHITECTURE BEHAV OF D2_4bit IS
BEGIN
--variable Enable:STD_LOGIC;
    PROCESS (VERT_SYNC)
    BEGIN
        IF RISING_EDGE(VERT_SYNC) THEN --add enable 
            IF SCORE_IN >= 0 AND SCORE_IN <= 9 THEN
                SCORE_OUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(SCORE_IN, 4));
		--Enable<='1;'
		--ELSE
		--Enable<='0';
            END IF;
        END IF;
--ENABLE_OUT<=ENABLE;
    END PROCESS;
END ARCHITECTURE BEHAV;

