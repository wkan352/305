library IEEE;
use  IEEE.STD_LOGIC_1164.all;
use  IEEE.STD_LOGIC_ARITH.all;
use  IEEE.STD_LOGIC_UNSIGNED.all;

entity text_display is
	port(	show_text : in std_logic;
	red_in, green_in, blue_in : in std_logic_vector(3 downto 0);
		pixel_row,pixel_col : in std_logic_vector(9 downto 0);
		red_out, green_out, blue_out : out std_logic_vector(3 downto 0));
end entity text_display;

architecture behav of text_display is

	type alphaArray is array (0 to 46, 0 to 314) of std_logic;
	signal welcome_alphaArray : alphaArray := (
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"111111111110000000000000001111111110000000000000000111111111111000001111111111111111111111111110000000011111111111000000000000000000000000000000000000000111111111111111110000000000000000000000000011111111111111110000000000000000000000011111111111110000000000000000000111111111111000000000011111111111111111111111111",
"111111111110000000000000001111111111000000000000001111111111111000001111111111111111111111111110000000011111111111000000000000000000000000000000000000111111111111111111111110000000000000000000011111111111111111111100000000000000000000011111111111110000000000000000001111111111111000000000011111111111111111111111111",
"111111111111000000000000001111111111000000000000001111111111111000001111111111111111111111111110000000011111111111000000000000000000000000000000000011111111111111111111111111100000000000000000111111111111111111111111000000000000000000011111111111110000000000000000001111111111111000000000011111111111111111111111111",
"111111111111000000000000001111111111000000000000001111111111110000001111111111111111111111111110000000011111111111000000000000000000000000000000001111111111111111111111111111110000000000000011111111111111111111111111100000000000000000011111111111111000000000000000011111111111111000000000011111111111111111111111111",
"111111111111000000000000011111111111000000000000001111111111110000001111111111111111111111111110000000011111111111000000000000000000000000000000011111111111111111111111111111110000000000000111111111111111111111111111111000000000000000011111111111111000000000000000011111111111111000000000011111111111111111111111111",
"111111111111000000000000011111111111100000000000011111111111110000001111111111111111111111111110000000011111111111000000000000000000000000000000111111111111111111111111111111100000000000001111111111111111111111111111111100000000000000011111111111111000000000000000011111111111111000000000011111111111111111111111111",
"111111111111100000000000011111111111100000000000011111111111100000001111111111111111111111111110000000011111111111000000000000000000000000000001111111111111111111111111111111100000000000011111111111111111111111111111111110000000000000011111111111111100000000000000111111111111111000000000011111111111111111111111111",
"011111111111100000000000011111111111100000000000011111111111100000001111111111111111111111111110000000011111111111000000000000000000000000000011111111111111111111111111111111000000000000111111111111111111111111111111111111000000000000011111111111111100000000000000111111111111111000000000011111111111111111111111111",
"011111111111100000000000111111111111100000000000011111111111100000001111111111111111111111111110000000011111111111000000000000000000000000000111111111111111111111111111111111000000000001111111111111111111111111111111111111000000000000011111111111111110000000000001111111111111111000000000011111111111111111111111111",
"011111111111100000000000111111111111110000000000111111111111100000001111111111111111111111111110000000011111111111000000000000000000000000001111111111111111111111111111111110000000000011111111111111111111111111111111111111100000000000011111111111111110000000000001111111111111111000000000011111111111111111111111111",
"011111111111110000000000111111111111110000000000111111111111000000001111111111100000000000000000000000011111111111000000000000000000000000011111111111111111111110011111111110000000000011111111111111111000001111111111111111110000000000011111111111111110000000000001111111111111111100000000011111111111000000000000000",
"001111111111110000000001111111111111110000000000111111111111000000001111111111100000000000000000000000011111111111000000000000000000000000011111111111111111000000000001111100000000000111111111111111100000000001111111111111110000000000111111111111111111000000000011111111111111111100000000011111111111000000000000000",
"001111111111110000000001111111111111111000000000111111111111000000001111111111100000000000000000000000011111111111000000000000000000000000111111111111111100000000000000001100000000000111111111111110000000000000111111111111111000000000111111111111111111000000000011111111111111111100000000011111111111000000000000000",
"001111111111110000000001111111111111111000000001111111111110000000001111111111100000000000000000000000011111111111000000000000000000000000111111111111111000000000000000000000000000001111111111111100000000000000011111111111111000000000111111111111111111100000000011111111111111111100000000011111111111000000000000000",
"000111111111111000000001111111111111111000000001111111111110000000001111111111100000000000000000000000011111111111000000000000000000000001111111111111110000000000000000000000000000001111111111111000000000000000001111111111111100000000111111111111111111100000000111111111111111111100000000011111111111000000000000000",
"000111111111111000000011111111111111111000000001111111111110000000001111111111100000000000000000000000011111111111000000000000000000000001111111111111100000000000000000000000000000011111111111111000000000000000000111111111111100000000111111111111111111100000000111111111111111111100000000011111111111000000000000000",
"000111111111111000000011111111111111111100000001111111111110000000001111111111100000000000000000000000011111111111000000000000000000000001111111111111000000000000000000000000000000011111111111110000000000000000000111111111111100000000111111111111111111110000001111111111111111111100000000011111111111000000000000000",
"000111111111111000000011111111111111111100000011111111111100000000001111111111100000000000000000000000011111111111000000000000000000000011111111111110000000000000000000000000000000011111111111110000000000000000000011111111111100000000111111111111111111110000001111111111111111111100000000011111111111000000000000000",
"000011111111111100000011111111111111111100000011111111111100000000001111111111111111111111111100000000011111111111000000000000000000000011111111111110000000000000000000000000000000011111111111100000000000000000000011111111111110000000111111111111111111110000001111111111111111111100000000011111111111111111111111111",
"000011111111111100000111111111111111111100000011111111111100000000001111111111111111111111111100000000011111111111000000000000000000000011111111111100000000000000000000000000000000011111111111100000000000000000000011111111111110000000111111111111111111111000011111111111111111111100000000011111111111111111111111111",
"000011111111111100000111111111111111111110000011111111111000000000001111111111111111111111111100000000011111111111000000000000000000000011111111111100000000000000000000000000000000111111111111100000000000000000000001111111111110000000111111111111111111111000011111111111111111111100000000011111111111111111111111111",
"000001111111111100000111111111111111111110000111111111111000000000001111111111111111111111111100000000011111111111000000000000000000000011111111111100000000000000000000000000000000111111111111100000000000000000000001111111111110000000111111111111111111111100111111111111111111111110000000011111111111111111111111111",
"000001111111111110000111111111111111111110000111111111111000000000001111111111111111111111111100000000011111111111000000000000000000000011111111111100000000000000000000000000000000111111111111100000000000000000000001111111111110000001111111111111111111111100111111111111111111111110000000011111111111111111111111111",
"000001111111111110001111111111111111111110000111111111111000000000001111111111111111111111111100000000011111111111000000000000000000000011111111111100000000000000000000000000000000111111111111000000000000000000000001111111111110000001111111111110111111111100111111111110111111111110000000011111111111111111111111111",
"000001111111111110001111111111011111111111000111111111110000000000001111111111111111111111111100000000011111111111000000000000000000000011111111111100000000000000000000000000000000111111111111000000000000000000000001111111111110000001111111111100111111111111111111111100111111111110000000011111111111111111111111111",
"000000111111111110001111111111001111111111001111111111110000000000001111111111111111111111111100000000011111111111000000000000000000000011111111111100000000000000000000000000000000111111111111100000000000000000000001111111111110000001111111111100111111111111111111111100111111111110000000011111111111111111111111111",
"000000111111111111001111111111001111111111001111111111110000000000001111111111111111111111111100000000011111111111000000000000000000000011111111111100000000000000000000000000000000111111111111100000000000000000000011111111111110000001111111111100011111111111111111111000111111111110000000011111111111111111111111111",
"000000111111111111011111111110001111111111101111111111100000000000001111111111111111111111111100000000011111111111000000000000000000000011111111111110000000000000000000000000000000011111111111100000000000000000000011111111111110000001111111111100011111111111111111111000111111111110000000011111111111111111111111111",
"000000011111111111011111111110000111111111101111111111100000000000001111111111100000000000000000000000011111111111000000000000000000000011111111111110000000000000000000000000000000011111111111100000000000000000000011111111111110000001111111111100011111111111111111111000111111111110000000011111111111000000000000000",
"000000011111111111011111111110000111111111111111111111100000000000001111111111100000000000000000000000011111111111000000000000000000000011111111111111000000000000000000000000000000011111111111110000000000000000000011111111111100000001111111111100001111111111111111110000111111111110000000011111111111000000000000000",
"000000011111111111111111111110000111111111111111111111100000000000001111111111100000000000000000000000011111111111000000000000000000000001111111111111000000000000000000000000000000011111111111110000000000000000000111111111111100000001111111111100001111111111111111110000111111111110000000011111111111000000000000000",
"000000011111111111111111111100000111111111111111111111000000000000001111111111100000000000000000000000011111111111000000000000000000000001111111111111100000000000000000000000000000011111111111111000000000000000001111111111111100000001111111111100001111111111111111110000111111111110000000011111111111000000000000000",
"000000001111111111111111111100000011111111111111111111000000000000001111111111100000000000000000000000011111111111000000000000000000000001111111111111110000000000000000000000000000001111111111111000000000000000001111111111111000000001111111111100000111111111111111100000111111111110000000011111111111000000000000000",
"000000001111111111111111111100000011111111111111111111000000000000001111111111100000000000000000000000011111111111000000000000000000000000111111111111111000000000000000001100000000001111111111111100000000000000011111111111111000000011111111111100000111111111111111100000111111111111000000011111111111000000000000000",
"000000001111111111111111111000000011111111111111111110000000000000001111111111100000000000000000000000011111111111000000000000000000000000111111111111111110000000000000011100000000000111111111111111000000000000111111111111111000000011111111111100000111111111111111100000111111111111000000011111111111000000000000000",
"000000000111111111111111111000000001111111111111111110000000000000001111111111100000000000000000000000011111111111000000000000000000000000011111111111111111100000000011111110000000000111111111111111110000000011111111111111110000000011111111111100000011111111111111000000111111111111000000011111111111000000000000000",
"000000000111111111111111111000000001111111111111111110000000000000001111111111111111111111111110000000011111111111111111111111111100000000001111111111111111111111111111111110000000000011111111111111111111111111111111111111110000000011111111111100000011111111111111000000011111111111000000011111111111111111111111111",
"000000000111111111111111111000000001111111111111111110000000000000001111111111111111111111111110000000011111111111111111111111111100000000001111111111111111111111111111111111000000000011111111111111111111111111111111111111100000000011111111111000000011111111111111000000011111111111000000011111111111111111111111111",
"000000000111111111111111110000000001111111111111111100000000000000001111111111111111111111111110000000011111111111111111111111111100000000000111111111111111111111111111111111000000000001111111111111111111111111111111111111000000000011111111111000000001111111111110000000011111111111000000011111111111111111111111111",
"000000000011111111111111110000000000111111111111111100000000000000001111111111111111111111111110000000011111111111111111111111111100000000000011111111111111111111111111111111100000000000111111111111111111111111111111111110000000000011111111111000000001111111111110000000011111111111000000011111111111111111111111111",
"000000000011111111111111110000000000111111111111111100000000000000001111111111111111111111111110000000011111111111111111111111111100000000000001111111111111111111111111111111100000000000011111111111111111111111111111111100000000000011111111111000000000111111111110000000011111111111000000011111111111111111111111111",
"000000000011111111111111100000000000111111111111111000000000000000001111111111111111111111111110000000011111111111111111111111111100000000000000111111111111111111111111111111110000000000001111111111111111111111111111111000000000000011111111111000000000111111111100000000011111111111000000011111111111111111111111111",
"000000000001111111111111100000000000011111111111111000000000000000001111111111111111111111111110000000011111111111111111111111111100000000000000001111111111111111111111111111110000000000000111111111111111111111111111110000000000000011111111111000000000111111111100000000011111111111000000011111111111111111111111111",
"000000000001111111111111100000000000011111111111111000000000000000001111111111111111111111111110000000011111111111111111111111111100000000000000000111111111111111111111111111100000000000000011111111111111111111111111100000000000000011111111111000000000011111111100000000011111111111000000011111111111111111111111111",
"000000000001111111111111100000000000011111111111111000000000000000001111111111111111111111111110000000011111111111111111111111111100000000000000000001111111111111111111111111000000000000000000111111111111111111111110000000000000000111111111111000000000011111111000000000011111111111100000011111111111111111111111111",
"000000000001111111111111000000000000011111111111110000000000000000001111111111111111111111111110000000011111111111111111111111111100000000000000000000011111111111111111111000000000000000000000001111111111111111111000000000000000000111111111111000000000011111111000000000011111111111100000011111111111111111111111111");

	
	Constant text_start_X: std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(162, 10);
	Constant text_end_X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(477, 10);
	
	Constant text_start_Y: std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(215, 10);
	Constant text_end_Y: std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(261, 10);	
	signal is_text : boolean;
	
begin
	is_text <= ((pixel_row >= text_start_Y) and (pixel_row < text_end_Y) and
			(pixel_col >= text_start_X) and (pixel_col < text_end_X) and 
			(welcome_alphaArray(CONV_INTEGER(unsigned(pixel_row - text_start_Y)) , CONV_INTEGER(unsigned(pixel_col - text_start_X))) = '1') and show_text = '1');
	
	red_out <= "1111" when (is_text =true) else red_in;
	green_out <= "1111" when (is_text =true) else green_in;
	blue_out <= "1111" when (is_text =true) else blue_in;
	
end architecture behav;