LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BIRD IS
	PORT (	LEFT_MOUSE, VERT_SYNC : IN STD_LOGIC;
		RED_IN, GREEN_IN, BLUE_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		PIXEL_ROW, PIXEL_COL : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		RED,GREEN,BLUE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ENTITY BIRD;

ARCHITECTURE BEHAV OF BIRD IS

	SIGNAL IS_BIRD : STD_LOGIC;
	CONSTANT BIRD_SIZE : INTEGER := 20;
	CONSTANT BIRD_X : INTEGER := 100;
	SIGNAL BIRD_Y : INTEGER := 239;
	
	SIGNAL ROW_INT : INTEGER;
	SIGNAL COL_INT : INTEGER;

BEGIN
	-- CONVERSIONS
	ROW_INT <= TO_INTEGER(UNSIGNED(PIXEL_ROW));
	COL_INT <= TO_INTEGER(UNSIGNED(PIXEL_COL)); 
	

	IS_BIRD <= '1' WHEN ( (ROW_INT >= BIRD_Y) AND (ROW_INT <= BIRD_Y + BIRD_SIZE) AND
			(COL_INT <= BIRD_X) AND (COL_INT >= BIRD_X - BIRD_SIZE) ) ELSE '0' ;
	
	RED <= "1111" WHEN IS_BIRD = '1' ELSE RED_IN;
	GREEN <= "1111" WHEN IS_BIRD ='1' ELSE GREEN_IN;
	BLUE <= "0000" WHEN IS_BIRD = '1' ELSE BLUE_IN;

	MOVE_BIRD: PROCESS(VERT_SYNC)
		VARIABLE CLICKED_ALREADY : STD_LOGIC := '0';
		VARIABLE GRAVITY : INTEGER := 0;
		VARIABLE BIRD_MOTION : INTEGER := 0;
		
	BEGIN
		IF(RISING_EDGE(VERT_SYNC)) THEN
			IF(LEFT_MOUSE ='1' AND CLICKED_ALREADY = '0') THEN
				BIRD_MOTION := -12;
				GRAVITY := 1;
				
			ELSE
				BIRD_MOTION := BIRD_MOTION + GRAVITY;
				
			END IF;
			
			IF((BIRD_Y <= (40 + BIRD_MOTION)) OR (BIRD_Y >= (438 - BIRD_SIZE))) THEN
				BIRD_Y <= 239;
				BIRD_MOTION := 0;
				GRAVITY := 0;
			ELSE
				BIRD_Y <= BIRD_Y + BIRD_MOTION;
			END IF;

			IF LEFT_MOUSE ='1' THEN
				CLICKED_ALREADY :='1';
				
			ELSE
				CLICKED_ALREADY := '0';
				
			END IF;
		END IF;
	END PROCESS MOVE_BIRD;
END ARCHITECTURE BEHAV;