LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BIRD IS
	PORT (	RED_IN, GREEN_IN, BLUE_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		BIRD_X, BIRD_Y : IN INTEGER;
		PIXEL_ROW, PIXEL_COL : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		RED,GREEN,BLUE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ENTITY BIRD;

ARCHITECTURE BEHAV OF BIRD IS

	SIGNAL IS_BIRD : STD_LOGIC;
	CONSTANT BIRD_SIZE : INTEGER := 20;
	
	SIGNAL ROW_INT : INTEGER;
	SIGNAL COL_INT : INTEGER;

BEGIN
	-- CONVERSIONS
	ROW_INT <= TO_INTEGER(UNSIGNED(PIXEL_ROW));
	COL_INT <= TO_INTEGER(UNSIGNED(PIXEL_COL)); 
	

	IS_BIRD <= '1' WHEN ( (ROW_INT >= BIRD_Y) AND (ROW_INT <= BIRD_Y + BIRD_SIZE) AND
			(COL_INT <= BIRD_X) AND (COL_INT >= BIRD_X - BIRD_SIZE) ) ELSE '0' ;
	
	RED <= "1111" WHEN IS_BIRD = '1' ELSE RED_IN;
	GREEN <= "1111" WHEN IS_BIRD ='1' ELSE GREEN_IN;
	BLUE <= "0000" WHEN IS_BIRD = '1' ELSE BLUE_IN;

END ARCHITECTURE BEHAV;

